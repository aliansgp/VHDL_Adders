
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity carry_generator is
	Port ( G : in  STD_LOGIC_VECTOR(15 downto 0);
			  P : in  STD_LOGIC_VECTOR(15 downto 0);
			  cin : STD_LOGIC;
           c : out  STD_LOGIC_VECTOR(15 downto 0));
end carry_generator;

architecture Behavioral of carry_generator is

begin
c(0) <= G(0) or (cin and P(0));
c(1) <= G(1) or (G(0) and P(1)) or (cin and P(0) and P(1));
c(2) <= G(2) or (G(1) and P(2)) or (G(0) and P(1) and P(2)) or (cin and P(0) and P(1) and P(2));
c(3) <= G(3) or (G(2) and P(3)) or (G(1) and P(2) and P(3)) or (G(0) and P(1) and P(2) and P(3)) or (cin and P(0) and P(1) and P(2) and P(3));
c(4) <= G(4) or (G(3) and P(4)) or (G(2) and P(3) and P(4)) or (G(1) and P(2) and P(3) and P(4)) or (p(0) and P(1) and P(2) and P(3) and P(4)) or (cin and p(0) and P(1) and P(2) and P(3) and P(4));
c(5) <= G(5) or (G(4) and P(5)) or (G(3) and P(4) and P(5)) or (G(2) and P(3) and P(4) and P(5)) or (p(1) and P(2) and P(3) and P(4) and P(5)) or (p(0) and p(1) and P(2) and P(3) and P(4) and P(5)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5));
c(6) <= G(6) or (G(5) and P(6)) or (G(4) and P(5) and P(6)) or (G(3) and P(4) and P(5) and P(6)) or (p(2) and P(3) and P(4) and P(5) and P(6)) or (p(1) and p(2) and P(3) and P(4) and P(5) and P(6)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6));
c(7) <= G(7) or (G(6) and P(7)) or (G(5) and P(6) and P(7)) or (G(4) and P(5) and P(6) and P(7)) or (p(3) and P(4) and P(5) and P(6) and P(7)) or (p(2) and p(3) and P(4) and P(5) and P(6) and P(7)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7));
c(8) <= G(8) or (G(7) and P(8)) or (G(6) and P(7) and P(8)) or (G(5) and P(6) and P(7) and P(8)) or (p(4) and P(5) and P(6) and P(7) and P(8)) or (p(3) and p(4) and P(5) and P(6) and P(7) and P(8)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8));
c(9) <= G(9) or (G(8) and P(9)) or (G(7) and P(8) and P(9)) or (G(6) and P(7) and P(8) and P(9)) or (p(5) and P(6) and P(7) and P(8) and P(9)) or (p(4) and p(5) and P(6) and P(7) and P(8) and P(9)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9));
c(10) <= G(10) or (G(9) and P(10)) or (G(8) and P(9) and P(10)) or (G(7) and P(8) and P(9) and P(10)) or (p(6) and P(7) and P(8) and P(9) and P(10)) or (p(5) and p(6) and P(7) and P(8) and P(9) and P(10)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10));
c(11) <= G(11) or (G(10) and P(11)) or (G(9) and P(10) and P(11)) or (G(8) and P(9) and P(10) and P(11)) or (p(7) and P(8) and P(9) and P(10) and P(11)) or (p(6) and p(7) and P(8) and P(9) and P(10) and P(11)) or (P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11));
c(12) <= G(12) or (G(11) and P(12)) or (G(10) and P(11) and P(12)) or (G(9) and P(10) and P(11) and P(12)) or (p(8) and P(9) and P(10) and P(11) and P(12)) or (p(7) and p(8) and P(9) and P(10) and P(11) and P(12)) or (P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12));
c(13) <= G(13) or (G(12) and P(13)) or (G(11) and P(12) and P(13)) or (G(10) and P(11) and P(12) and P(13)) or (p(9) and P(10) and P(11) and P(12) and P(13)) or (p(8) and p(9) and P(10) and P(11) and P(12) and P(13)) or (P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(12) and P(13)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13));
c(14) <= G(14) or (G(13) and P(14)) or (G(12) and P(13) and P(14)) or (G(11) and P(12) and P(13) and P(14)) or (p(10) and P(11) and P(12) and P(13) and P(14)) or (p(9) and p(10) and P(11) and P(12) and P(13) and P(14)) or (P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14));
c(15) <= G(15) or (G(14) and P(15)) or (G(13) and P(14) and P(15)) or (G(12) and P(13) and P(14) and P(15)) or (p(11) and P(12) and P(13) and P(14) and P(15)) or (p(10) and p(11) and P(12) and P(13) and P(14) and P(15)) or (P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15)) or (cin and P(0) and P(1) and P(2) and P(3) and P(4) and P(5) and P(6) and P(7) and P(8) and P(9) and P(10) and P(11) and P(12) and P(13) and P(14) and P(15));
end Behavioral;

